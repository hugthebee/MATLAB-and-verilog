magic
tech scmos
timestamp 1669655132
<< nwell >>
rect -21 3 32 20
rect 40 3 93 20
<< ntransistor >>
rect -5 -33 -2 -28
rect 13 -33 16 -28
rect 63 -33 67 -28
<< ptransistor >>
rect -5 9 -2 14
rect 13 9 16 14
rect 63 9 67 14
<< ndiffusion >>
rect -10 -33 -5 -28
rect -2 -33 13 -28
rect 16 -33 20 -28
rect 51 -33 63 -28
rect 67 -33 81 -28
<< pdiffusion >>
rect -10 9 -5 14
rect -2 9 4 14
rect 9 9 13 14
rect 16 9 20 14
rect 51 9 63 14
rect 67 9 81 14
<< ndcontact >>
rect -15 -33 -10 -28
rect 20 -33 25 -28
rect 46 -33 51 -28
rect 81 -33 86 -28
<< pdcontact >>
rect -15 9 -10 14
rect 4 9 9 14
rect 20 9 25 14
rect 46 9 51 14
rect 81 9 86 14
<< psubstratepcontact >>
rect -10 -45 -3 -38
rect 9 -45 16 -38
rect 55 -45 62 -38
rect 74 -45 81 -38
<< nwsc >>
rect -10 26 -3 33
rect 7 26 14 33
rect 49 26 56 33
rect 73 26 80 33
<< polysilicon >>
rect -5 14 -2 25
rect 13 14 16 25
rect 63 14 67 24
rect -5 -28 -2 9
rect 13 -28 16 9
rect 63 -4 67 9
rect 30 -9 67 -4
rect 63 -28 67 -9
rect -5 -36 -2 -33
rect 13 -36 16 -33
rect 63 -36 67 -33
<< polycontact >>
rect 25 -9 30 -4
<< metal1 >>
rect -15 14 -10 33
rect -3 26 7 33
rect 14 26 49 33
rect 56 26 73 33
rect 80 26 93 33
rect 20 14 25 26
rect 46 14 51 26
rect 4 -4 9 9
rect 4 -9 25 -4
rect 20 -28 25 -9
rect 81 -28 86 9
rect -15 -45 -10 -33
rect 46 -38 51 -33
rect -3 -45 9 -38
rect 16 -45 55 -38
rect 62 -45 74 -38
rect 81 -45 86 -38
<< end >>
