magic
tech scmos
timestamp 1669654258
<< metal1 >>
rect -44 67 -5 71
rect -23 60 -7 64
rect 175 61 189 65
rect 12 -40 33 -36
rect 12 -47 33 -43
rect 125 -45 143 -40
use xor  xor_0
timestamp 1669650328
transform 1 0 3 0 1 37
box -21 -26 191 110
use and  and_0
timestamp 1669650498
transform 1 0 45 0 1 -68
box -27 -2 102 66
<< labels >>
rlabel space -38 60 -22 64 3 B
rlabel space -55 67 -41 71 3 A
rlabel space 189 61 203 65 7 SUM
rlabel space 128 -49 146 -44 1 CARRY
rlabel space 11 -43 20 -39 1 A
rlabel space 11 -50 20 -46 1 B
<< end >>
