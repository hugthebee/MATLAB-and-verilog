magic
tech scmos
timestamp 1669665579
<< nwell >>
rect -46 3 96 21
<< ntransistor >>
rect -28 -31 -25 -25
rect 3 -31 6 -25
rect 41 -31 45 -25
rect 73 -31 77 -25
<< ptransistor >>
rect -28 9 -24 15
rect 4 9 8 15
rect 41 9 45 15
rect 73 9 77 15
<< ndiffusion >>
rect -38 -26 -28 -25
rect -38 -30 -34 -26
rect -30 -30 -28 -26
rect -38 -31 -28 -30
rect -25 -26 -10 -25
rect -25 -30 -21 -26
rect -17 -30 -10 -26
rect -25 -31 -10 -30
rect -6 -26 3 -25
rect -6 -30 -4 -26
rect 0 -30 3 -26
rect -6 -31 3 -30
rect 6 -26 22 -25
rect 6 -30 15 -26
rect 19 -30 22 -26
rect 6 -31 22 -30
rect 27 -26 41 -25
rect 27 -30 29 -26
rect 33 -30 41 -26
rect 27 -31 41 -30
rect 45 -26 55 -25
rect 45 -30 49 -26
rect 53 -30 55 -26
rect 45 -31 55 -30
rect 63 -26 73 -25
rect 63 -30 65 -26
rect 69 -30 73 -26
rect 63 -31 73 -30
rect 77 -26 91 -25
rect 77 -30 84 -26
rect 88 -30 91 -26
rect 77 -31 91 -30
<< pdiffusion >>
rect -39 14 -28 15
rect -39 10 -34 14
rect -30 10 -28 14
rect -39 9 -28 10
rect -24 14 -11 15
rect -24 10 -21 14
rect -17 10 -11 14
rect -24 9 -11 10
rect -7 14 4 15
rect -7 10 -4 14
rect 0 10 4 14
rect -7 9 4 10
rect 8 14 21 15
rect 8 10 15 14
rect 19 10 21 14
rect 8 9 21 10
rect 27 14 41 15
rect 27 10 29 14
rect 33 10 41 14
rect 27 9 41 10
rect 45 14 55 15
rect 45 10 49 14
rect 53 10 55 14
rect 45 9 55 10
rect 62 14 73 15
rect 62 10 65 14
rect 69 10 73 14
rect 62 9 73 10
rect 77 14 90 15
rect 77 10 84 14
rect 88 10 90 14
rect 77 9 90 10
<< ndcontact >>
rect -34 -30 -30 -26
rect -21 -30 -17 -26
rect -4 -30 0 -26
rect 15 -30 19 -26
rect 29 -30 33 -26
rect 49 -30 53 -26
rect 65 -30 69 -26
rect 84 -30 88 -26
<< pdcontact >>
rect -34 10 -30 14
rect -21 10 -17 14
rect -4 10 0 14
rect 15 10 19 14
rect 29 10 33 14
rect 49 10 53 14
rect 65 10 69 14
rect 84 10 88 14
<< psubstratepcontact >>
rect 36 -48 40 -44
rect 58 -48 62 -44
<< nwsc >>
rect 40 24 46 30
rect 58 24 64 30
<< polysilicon >>
rect -58 31 8 34
rect -58 -39 -55 31
rect -28 15 -24 23
rect 4 15 8 31
rect 41 15 45 22
rect 73 15 77 23
rect -28 -16 -24 9
rect 4 0 8 9
rect -28 -19 6 -16
rect -28 -25 -25 -22
rect 3 -25 6 -19
rect 41 -25 45 9
rect 73 -8 77 9
rect 67 -15 77 -8
rect 73 -25 77 -15
rect -28 -39 -25 -31
rect -58 -42 -25 -39
rect -28 -67 -25 -42
rect 3 -55 6 -31
rect 41 -36 45 -31
rect 73 -55 77 -31
rect 3 -58 77 -55
rect 105 -67 114 -8
rect -28 -70 114 -67
<< polycontact >>
rect 35 -14 41 -8
rect 99 -15 105 -8
<< metal1 >>
rect -34 36 26 40
rect -34 14 -30 36
rect -34 -26 -30 10
rect -21 24 19 29
rect -21 14 -17 24
rect 15 14 19 24
rect -21 -26 -17 10
rect -4 -26 0 10
rect 23 -8 26 36
rect 29 24 40 30
rect 46 24 58 30
rect 64 24 69 30
rect 29 14 33 24
rect 65 14 69 24
rect 23 -14 35 -8
rect 49 -19 53 10
rect 23 -23 53 -19
rect -4 -38 0 -30
rect 23 -38 26 -23
rect 49 -26 53 -23
rect 84 -8 88 10
rect 84 -15 99 -8
rect 84 -26 88 -15
rect -4 -42 26 -38
rect 29 -44 33 -30
rect 65 -44 69 -30
rect 29 -48 36 -44
rect 40 -48 58 -44
rect 62 -48 69 -44
<< end >>
