magic
tech scmos
timestamp 1669666639
<< error_s >>
rect 609 483 631 484
rect 615 477 628 479
rect 813 443 817 444
rect 821 443 837 444
rect 819 437 834 439
rect 819 436 821 437
rect 822 434 824 436
rect 1306 421 1328 422
rect 1312 415 1325 417
rect 1510 381 1514 382
rect 1518 381 1534 382
rect 1516 375 1531 377
rect 1516 374 1518 375
rect 1519 372 1521 374
rect 845 337 852 340
rect 862 337 869 340
rect 904 337 911 340
rect 928 337 935 340
rect 948 335 949 336
rect 1240 306 1241 311
rect 1240 299 1242 306
rect 1542 275 1549 278
rect 1559 275 1566 278
rect 1601 275 1608 278
rect 1625 275 1632 278
rect 1645 273 1646 274
rect 845 262 851 265
rect 864 262 868 265
rect 910 262 916 269
rect 929 262 934 265
rect 947 260 948 261
rect 839 253 841 260
rect 1542 200 1548 203
rect 1561 200 1565 203
rect 1607 200 1613 207
rect 1626 200 1631 203
rect 318 199 343 200
rect 1644 198 1645 199
rect 324 193 340 195
rect 1536 191 1538 198
rect 1989 157 2014 158
rect 1995 151 2011 153
rect 699 150 721 151
rect 705 144 718 146
rect 903 110 907 111
rect 911 110 927 111
rect 909 104 924 106
rect 725 72 755 74
rect 899 44 901 104
rect 909 103 911 104
rect 912 101 914 103
rect 1336 102 1358 103
rect 1342 96 1355 98
rect 1540 62 1544 63
rect 1548 62 1564 63
rect 1546 56 1561 58
rect 1546 55 1548 56
rect 1549 53 1551 55
rect 1395 18 1426 19
rect 1431 18 1435 19
rect 935 4 942 7
rect 952 4 959 7
rect 994 4 1001 7
rect 1018 4 1025 7
rect 1038 2 1039 3
rect -17 -17 -7 -12
rect -4 -17 11 -12
rect 18 -17 23 -16
rect 44 -17 61 -12
rect 65 -17 84 -12
rect -17 -31 -16 -17
rect -12 -21 -5 -19
rect 5 -21 12 -19
rect 47 -21 54 -19
rect 71 -21 78 -19
rect -12 -26 -5 -22
rect 7 -26 12 -22
rect 53 -26 54 -22
rect 72 -26 78 -22
rect -7 -29 -5 -27
rect 11 -29 14 -27
rect 138 -37 145 -36
rect 157 -37 164 -36
rect 203 -37 210 -36
rect 222 -37 229 -36
rect 133 -54 135 -42
rect 1572 -44 1579 -41
rect 1589 -44 1596 -41
rect 1631 -44 1638 -41
rect 1655 -44 1662 -41
rect 1675 -46 1676 -45
rect 316 -50 341 -49
rect 322 -56 338 -54
rect 704 -59 705 -47
rect 935 -71 941 -68
rect 954 -71 958 -68
rect 1000 -71 1006 -64
rect 1019 -71 1024 -68
rect 1037 -73 1038 -72
rect 929 -80 931 -73
rect 1985 -74 2007 -73
rect 1991 -80 2004 -78
rect -17 -85 -7 -80
rect -4 -85 11 -80
rect 18 -85 23 -84
rect 44 -85 61 -80
rect 65 -85 84 -80
rect 152 -84 168 -82
rect 173 -84 178 -82
rect -12 -89 -5 -87
rect 5 -89 12 -87
rect 47 -89 54 -87
rect 71 -89 78 -87
rect -12 -94 -5 -90
rect 7 -94 12 -90
rect 53 -94 54 -90
rect 72 -94 78 -90
rect -7 -97 -5 -95
rect 11 -97 14 -95
rect 86 -97 87 -94
rect 701 -107 712 -105
rect 762 -107 773 -105
rect 1572 -119 1578 -116
rect 1591 -119 1595 -116
rect 1637 -119 1643 -112
rect 2206 -114 2213 -113
rect 1656 -119 1661 -116
rect 2195 -119 2210 -118
rect 1674 -121 1675 -120
rect 1566 -128 1568 -121
rect 133 -140 135 -128
rect 1301 -131 1357 -129
rect 1362 -131 1400 -129
rect -17 -153 -7 -148
rect -4 -153 11 -148
rect 18 -153 23 -152
rect 44 -153 61 -148
rect 65 -153 84 -148
rect -17 -167 -15 -153
rect -12 -157 -5 -155
rect 5 -157 12 -155
rect 47 -157 54 -155
rect 71 -157 78 -155
rect -12 -162 -5 -158
rect 7 -162 12 -158
rect 53 -162 54 -158
rect 72 -162 78 -158
rect -7 -165 -5 -163
rect 11 -165 14 -163
rect 152 -170 168 -168
rect 173 -170 178 -168
rect 2185 -180 2187 -119
rect 2195 -121 2197 -119
rect 2202 -120 2210 -119
rect 2198 -123 2200 -121
rect 133 -229 135 -217
rect 2221 -220 2228 -217
rect 2238 -220 2245 -217
rect 2280 -220 2287 -217
rect 2304 -220 2311 -217
rect 2324 -222 2325 -221
rect 1418 -281 1440 -280
rect 319 -284 344 -283
rect 1424 -287 1437 -285
rect 325 -290 341 -288
rect 2221 -295 2227 -292
rect 2240 -295 2244 -292
rect 2286 -295 2292 -288
rect 2305 -295 2310 -292
rect 2323 -297 2324 -296
rect 2215 -304 2217 -297
rect 1622 -321 1626 -320
rect 1630 -321 1646 -320
rect 1628 -327 1643 -325
rect 1628 -328 1630 -327
rect 1631 -330 1633 -328
rect 1444 -359 1474 -357
rect 777 -427 799 -426
rect 1654 -427 1661 -424
rect 1671 -427 1678 -424
rect 1713 -427 1720 -424
rect 1737 -427 1744 -424
rect 1757 -429 1758 -428
rect 783 -433 796 -431
rect 773 -444 775 -441
rect 991 -467 1005 -466
rect 987 -473 1002 -471
rect 987 -474 989 -473
rect 990 -476 992 -474
rect 1418 -495 1419 -483
rect 1654 -502 1660 -499
rect 1673 -502 1677 -499
rect 1719 -502 1725 -495
rect 2000 -498 2022 -497
rect 1738 -502 1743 -499
rect 1756 -504 1757 -503
rect 2006 -504 2019 -502
rect 803 -505 833 -504
rect 1648 -511 1650 -504
rect 2204 -538 2208 -536
rect 2212 -538 2217 -536
rect 2221 -538 2228 -537
rect 2210 -543 2225 -542
rect 2210 -545 2212 -543
rect 2217 -544 2225 -543
rect 2213 -547 2215 -545
rect 1013 -573 1020 -570
rect 1030 -573 1037 -570
rect 1072 -573 1079 -570
rect 1096 -573 1103 -570
rect 1116 -575 1117 -574
rect 608 -613 610 -606
rect 1013 -648 1019 -645
rect 1032 -648 1036 -645
rect 1078 -648 1084 -641
rect 2236 -644 2243 -641
rect 2253 -644 2260 -641
rect 2295 -644 2302 -641
rect 2319 -644 2326 -641
rect 1097 -648 1102 -645
rect 2339 -646 2340 -645
rect 1115 -650 1116 -649
rect 1007 -657 1009 -650
rect 1779 -689 1780 -677
rect 2236 -719 2242 -716
rect 2255 -719 2259 -716
rect 2301 -719 2307 -712
rect 2320 -719 2325 -716
rect 2338 -721 2339 -720
rect 2230 -728 2232 -721
<< metal1 >>
rect 568 477 588 481
rect 568 422 572 477
rect 585 470 611 474
rect 585 422 590 470
rect 781 437 831 441
rect 568 418 637 422
rect 585 411 590 418
rect 585 406 623 411
rect 514 350 522 354
rect 514 343 522 347
rect 618 345 623 406
rect 633 350 637 418
rect 626 345 678 350
rect 633 255 637 345
rect 673 264 678 345
rect 781 330 785 437
rect 1032 431 1044 435
rect 1272 414 1286 419
rect 1209 406 1229 410
rect 770 326 820 330
rect 770 264 774 326
rect 1209 270 1213 406
rect 1225 401 1229 406
rect 1272 401 1277 414
rect 1302 401 1306 411
rect 1225 397 1306 401
rect 1272 357 1277 397
rect 1494 375 1524 379
rect 1272 352 1345 357
rect 1228 306 1238 310
rect 1340 306 1345 352
rect 1229 299 1239 303
rect 1340 301 1346 306
rect 1341 270 1346 301
rect 1494 270 1498 375
rect 1728 369 1755 373
rect 1062 266 1516 270
rect 673 260 811 264
rect 770 255 774 260
rect 601 251 811 255
rect 267 193 302 197
rect 267 106 271 193
rect 111 102 271 106
rect 279 186 323 190
rect 529 187 542 191
rect -34 44 -20 48
rect -34 37 -20 41
rect 87 39 100 44
rect 111 0 116 102
rect 279 90 284 186
rect 279 86 359 90
rect 125 36 133 40
rect 279 36 284 86
rect 601 85 605 251
rect 770 238 774 251
rect 617 234 775 238
rect 617 85 621 234
rect 1209 192 1213 266
rect 1341 203 1346 266
rect 1759 204 1948 208
rect 1341 198 1506 203
rect 1497 192 1505 195
rect 1155 191 1505 192
rect 1155 188 1501 191
rect 125 29 133 33
rect 238 31 284 36
rect 326 79 357 83
rect 482 81 621 85
rect 667 144 682 148
rect 326 0 329 79
rect 111 -3 329 0
rect -33 -24 -19 -20
rect 111 -24 116 -3
rect 443 -4 450 13
rect -33 -31 -19 -27
rect 87 -29 116 -24
rect 121 -9 300 -6
rect 121 -34 124 -9
rect 114 -37 124 -34
rect 114 -85 119 -37
rect 124 -47 132 -43
rect 124 -54 132 -50
rect 236 -52 277 -47
rect 273 -59 277 -52
rect 297 -56 300 -9
rect 601 -59 605 81
rect 667 1 671 144
rect 692 71 696 141
rect 893 104 917 108
rect 692 66 850 71
rect 273 -63 321 -59
rect 525 -63 605 -59
rect 641 -1 671 1
rect 845 -1 850 66
rect 893 5 898 104
rect 1155 102 1159 188
rect 1944 155 1948 204
rect 1944 151 1979 155
rect 1944 147 1948 151
rect 1119 98 1159 102
rect 1874 143 1995 147
rect 2205 145 2223 149
rect 1256 96 1319 100
rect 1256 16 1260 96
rect 1331 92 1333 93
rect 1311 87 1335 92
rect 1311 32 1316 87
rect 1501 56 1557 60
rect 1311 27 1431 32
rect 1426 16 1431 27
rect 1501 16 1505 56
rect 1874 54 1878 143
rect 1757 50 1878 54
rect 1874 41 1878 50
rect 1944 48 1948 143
rect 1944 44 2032 48
rect 1874 37 2037 41
rect 2154 39 2206 44
rect 1189 12 1505 16
rect 893 2 929 5
rect 641 -4 910 -1
rect -31 -92 -17 -88
rect 114 -89 268 -85
rect 114 -92 119 -89
rect -31 -99 -17 -95
rect 86 -97 119 -92
rect 127 -95 257 -92
rect 127 -105 130 -95
rect 107 -108 130 -105
rect -32 -160 -18 -156
rect 107 -160 110 -108
rect 253 -119 257 -95
rect 265 -103 268 -89
rect 273 -94 277 -63
rect 273 -97 325 -94
rect 265 -106 317 -103
rect 253 -123 308 -119
rect 124 -133 132 -129
rect 124 -140 132 -136
rect 236 -138 292 -133
rect -32 -167 -18 -163
rect 87 -165 110 -160
rect 107 -171 110 -165
rect 107 -175 282 -171
rect 124 -222 132 -218
rect 124 -229 132 -225
rect 234 -541 239 -222
rect 277 -400 282 -175
rect 287 -293 292 -138
rect 304 -289 308 -123
rect 314 -166 317 -106
rect 322 -159 325 -97
rect 322 -163 369 -159
rect 641 -163 646 -4
rect 314 -170 356 -166
rect 481 -168 646 -163
rect 667 -103 671 -4
rect 694 -52 702 -48
rect 845 -52 850 -4
rect 879 -5 910 -4
rect 694 -59 702 -55
rect 805 -57 898 -52
rect 893 -73 898 -57
rect 1189 -63 1193 12
rect 1151 -67 1193 -63
rect 893 -103 897 -76
rect 667 -107 897 -103
rect 667 -292 671 -107
rect 1256 -127 1260 12
rect 1285 -66 1296 -62
rect 1426 -66 1431 12
rect 1501 -49 1505 12
rect 1501 -53 1544 -49
rect 1285 -73 1296 -69
rect 1397 -71 1463 -66
rect 1458 -116 1463 -71
rect 1927 -80 1968 -76
rect 1927 -111 1931 -80
rect 1789 -115 1931 -111
rect 1960 -88 1985 -84
rect 1458 -121 1544 -116
rect 1227 -131 1538 -127
rect 833 -234 841 -230
rect 833 -241 841 -237
rect 945 -239 1128 -234
rect 287 -297 329 -293
rect 531 -296 671 -292
rect 287 -393 292 -297
rect 1123 -298 1128 -239
rect 1227 -298 1231 -131
rect 1393 -298 1398 -283
rect 1413 -298 1418 -291
rect 1926 -292 1930 -115
rect 1960 -292 1964 -88
rect 2201 -114 2206 39
rect 2180 -119 2206 -114
rect 2181 -225 2184 -119
rect 2410 -126 2428 -122
rect 2181 -228 2199 -225
rect 1926 -296 2187 -292
rect 1123 -303 1418 -298
rect 1960 -300 1964 -296
rect 287 -397 358 -393
rect 277 -404 358 -400
rect 484 -402 563 -397
rect 558 -507 563 -402
rect 631 -431 760 -428
rect 631 -507 636 -431
rect 768 -440 777 -436
rect 709 -441 775 -440
rect 709 -444 772 -441
rect 709 -507 714 -444
rect 965 -473 1001 -470
rect 965 -507 970 -473
rect 1227 -475 1231 -303
rect 1344 -422 1349 -303
rect 1393 -360 1398 -303
rect 1960 -304 2190 -300
rect 1603 -327 1637 -323
rect 1603 -360 1607 -327
rect 1960 -329 1964 -304
rect 1838 -333 1964 -329
rect 1368 -364 1607 -360
rect 1368 -422 1372 -364
rect 1393 -390 1398 -364
rect 1393 -395 1547 -390
rect 1542 -422 1547 -395
rect 1344 -427 1584 -422
rect 1198 -479 1231 -475
rect 558 -512 970 -507
rect 631 -541 636 -512
rect 709 -541 714 -512
rect 234 -546 782 -541
rect 597 -606 605 -602
rect 709 -606 714 -546
rect 777 -606 782 -546
rect 963 -578 968 -512
rect 963 -583 987 -578
rect 597 -613 607 -609
rect 709 -611 966 -606
rect 777 -657 782 -611
rect 962 -647 965 -611
rect 1368 -640 1372 -427
rect 1406 -488 1416 -484
rect 1542 -488 1547 -427
rect 1406 -495 1416 -491
rect 1516 -493 1547 -488
rect 1542 -506 1547 -493
rect 1579 -499 1584 -427
rect 1603 -432 1607 -364
rect 2438 -401 2442 -287
rect 2217 -405 2442 -401
rect 1603 -436 1628 -432
rect 1870 -498 1973 -494
rect 1579 -500 1593 -499
rect 1969 -500 1973 -498
rect 1579 -503 1618 -500
rect 1969 -504 1980 -500
rect 1542 -507 1604 -506
rect 1542 -511 1619 -507
rect 1230 -644 1372 -640
rect 962 -650 980 -647
rect 970 -657 976 -654
rect 778 -660 973 -657
rect 1768 -682 1777 -678
rect 1975 -682 1979 -504
rect 1993 -682 1998 -507
rect 2217 -539 2221 -405
rect 2182 -543 2221 -539
rect 2183 -649 2186 -543
rect 2424 -550 2451 -546
rect 2183 -652 2207 -649
rect 1768 -689 1777 -685
rect 1880 -687 1998 -682
rect 1975 -717 1979 -687
rect 1993 -717 1998 -687
rect 2457 -715 2483 -711
rect 1975 -721 2203 -717
rect 1993 -729 1998 -721
rect 2197 -729 2202 -725
rect 1993 -734 2202 -729
use and  and_8
timestamp 1669655132
transform 1 0 540 0 1 322
box -21 -45 93 33
use and  and_0
timestamp 1669655132
transform 1 0 -2 0 1 16
box -21 -45 93 33
use and  and_4
timestamp 1669655132
transform 1 0 148 0 1 8
box -21 -45 93 33
use ha  ha_1
timestamp 1669666639
transform 1 0 345 0 1 126
box -55 -113 203 77
use fa  fa_0
timestamp 1669666639
transform 1 0 968 0 1 292
box -387 -105 111 195
use and  and_12
timestamp 1669655132
transform 1 0 1255 0 1 278
box -21 -45 93 33
use and  and_1
timestamp 1669655132
transform 1 0 -2 0 1 -52
box -21 -45 93 33
use and  and_5
timestamp 1669655132
transform 1 0 148 0 1 -75
box -21 -45 93 33
use and  and_2
timestamp 1669655132
transform 1 0 -2 0 1 -120
box -21 -45 93 33
use and  and_3
timestamp 1669655132
transform 1 0 -2 0 1 -188
box -21 -45 93 33
use and  and_6
timestamp 1669655132
transform 1 0 148 0 1 -161
box -21 -45 93 33
use and  and_7
timestamp 1669655132
transform 1 0 148 0 1 -250
box -21 -45 93 33
use ha  ha_0
timestamp 1669666639
transform 1 0 343 0 1 -123
box -55 -113 203 77
use fa  fa_3
timestamp 1669666639
transform 1 0 1665 0 1 230
box -387 -105 111 195
use and  and_9
timestamp 1669655132
transform 1 0 719 0 1 -80
box -21 -45 93 33
use ha  ha_3
timestamp 1669666639
transform 1 0 2016 0 1 84
box -55 -113 203 77
use fa  fa_1
timestamp 1669666639
transform 1 0 1058 0 1 -41
box -387 -105 111 195
use and  and_13
timestamp 1669655132
transform 1 0 1311 0 1 -94
box -21 -45 93 33
use fa  fa_4
timestamp 1669666639
transform 1 0 1695 0 1 -89
box -387 -105 111 195
use ha  ha_2
timestamp 1669666639
transform 1 0 346 0 1 -357
box -55 -113 203 77
use and  and_11
timestamp 1669655132
transform 1 0 859 0 1 -262
box -21 -45 93 33
use and  and_10
timestamp 1669655132
transform 1 0 623 0 1 -634
box -21 -45 93 33
use fa  fa_2
timestamp 1669666639
transform 1 0 1136 0 1 -618
box -387 -105 111 195
use fa  fa_6
timestamp 1669666639
transform 1 0 2344 0 1 -265
box -387 -105 111 195
use and  and_14
timestamp 1669655132
transform 1 0 1433 0 1 -516
box -21 -45 93 33
use fa  fa_5
timestamp 1669666639
transform 1 0 1777 0 1 -472
box -387 -105 111 195
use and  and_15
timestamp 1669655132
transform 1 0 1794 0 1 -710
box -21 -45 93 33
use fa  fa_7
timestamp 1669666639
transform 1 0 2359 0 1 -689
box -387 -105 111 195
<< labels >>
rlabel space -44 44 -30 48 3 a0
rlabel space -34 34 -20 38 1 b0
rlabel space -33 -34 -19 -30 1 b0
rlabel space -35 -27 -21 -23 1 a1
rlabel space -35 -95 -21 -91 1 a2
rlabel space -35 -102 -21 -98 1 b0
rlabel space -33 -163 -19 -159 1 a3
rlabel space -32 -170 -18 -166 1 b0
rlabel space 90 35 103 40 1 p0
rlabel space 123 33 131 37 1 a0
rlabel space 125 26 133 30 1 b1
rlabel space 124 -50 132 -46 1 a1
rlabel space 124 -57 132 -53 1 b1
rlabel space 124 -136 132 -132 1 a2
rlabel space 123 -143 131 -139 1 b1
rlabel space 123 -225 131 -221 1 a3
rlabel space 123 -232 131 -228 1 b1
rlabel space 514 347 522 351 1 a0
rlabel space 514 340 522 344 1 b2
rlabel space 694 -55 702 -51 1 a1
rlabel space 694 -62 702 -58 1 b2
rlabel space 597 -609 605 -605 1 a2
rlabel space 597 -616 605 -612 1 b1
rlabel space 833 -237 841 -233 1 a3
rlabel space 834 -244 842 -240 1 b1
rlabel space 1034 428 1046 432 1 p2
rlabel space 1228 303 1238 307 1 a0
rlabel space 1229 296 1239 300 1 b3
rlabel space 1284 -69 1295 -65 1 a1
rlabel space 1284 -76 1295 -72 1 b3
rlabel space 1406 -490 1416 -486 1 a2
rlabel space 1406 -497 1416 -493 1 b3
rlabel space 1743 367 1755 370 1 p3
rlabel space 1768 -685 1777 -681 1 a3
rlabel space 1768 -692 1777 -688 1 b3
rlabel space 2214 142 2223 146 1 p4
rlabel space 2419 -129 2428 -125 1 p5
rlabel space 2442 -553 2451 -549 1 p6
rlabel space 2483 -715 2492 -711 7 p7
<< end >>
